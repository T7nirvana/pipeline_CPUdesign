`include "ctrl_encode_def.v"
module ID_EXT( Imm16, EXTOp, Imm32);
    
   input  [15:0] Imm16;
   input         EXTOp;
   output [31:0] Imm32;
   
   reg [31:0] Imm32;
    
   always @(*) begin
      case (EXTOp)
         `EXT_ZERO:    Imm32 = {16'd0, Imm16};
         `EXT_SIGNED:  Imm32 = {{16{Imm16[15]}}, Imm16};
         default: ;
      endcase
   end // end always
    
endmodule
